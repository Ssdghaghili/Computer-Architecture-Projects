module InstDataMemory (input clk,input reset,input [31:0] addr,data_in,input write_en,output reg[31:0] data_out);

  //dataMemory starts from mem[1024] to mem[4095]
//0000000 00010 00011 010 00111 0110011
  reg [7:0] mem [262143:0];
  assign data_out = {mem[addr+3],mem[addr+2],mem[addr+1],mem[addr]};

  always @(posedge clk) begin
    if (write_en)
    begin
      mem[addr] <= data_in[7:0];
      mem[addr+1] <= data_in[15:8];
      mem[addr+2] <= data_in[23:16];
      mem[addr+3] <= data_in[31:24];
    end
  end

  always @(reset)
    begin
        if(reset == 1)
        begin 

            // Setting arr = [12 , 1, -150 , 10 , 56 , 79 , 60 , 41 , 36 , 69] to memory using
            // addi x2 , zero , <number> and lw
            {mem[3],mem[2],mem[1],mem[0]} =32'b0000_0000_1100_00000_000_00010_0010011 ; 
            {mem[7],mem[6],mem[5],mem[4]} =32'b0100000_00010_00000_010_00000_0100011 ;//sw

            {mem[11],mem[10],mem[9],mem[8]} =32'b0000_0000_0001_00000_000_00010_0010011 ;
            {mem[15],mem[14],mem[13],mem[12]} =32'b0100000_00010_00000_010_00100_0100011 ;//sw

            {mem[19],mem[18],mem[17],mem[16]} =32'b1111_0110_1010_00000_000_00010_0010011 ;
            {mem[23],mem[22],mem[21],mem[20]} =32'b0100000_00010_00000_010_01000_0100011 ;//sw  

            {mem[27],mem[26],mem[25],mem[24]} =32'b0000_0000_1010_00000_000_00010_0010011 ;
            {mem[31],mem[30],mem[29],mem[28]} =32'b0100000_00010_00000_010_01100_0100011 ;//sw

            {mem[35],mem[34],mem[33],mem[32]} =32'b0000_0011_1000_00000_000_00010_0010011 ;
            {mem[39],mem[38],mem[37],mem[36]} =32'b0100000_00010_00000_010_10000_0100011 ;//sw

            {mem[43],mem[42],mem[41],mem[40]} =32'b0000_0100_1111_00000_000_00010_0010011 ;
            {mem[47],mem[46],mem[45],mem[44]} =32'b0100000_00010_00000_010_10100_0100011 ;//sw

            {mem[51],mem[50],mem[49],mem[48]} =32'b0000_0011_1100_00000_000_00010_0010011 ;
            {mem[55],mem[54],mem[53],mem[52]} =32'b0100000_00010_00000_010_11000_0100011 ;//sw

            {mem[59],mem[58],mem[57],mem[56]} =32'b0000_0010_1001_00000_000_00010_0010011 ;
            {mem[63],mem[62],mem[61],mem[60]} =32'b0100000_00010_00000_010_11100_0100011 ;//sw

            {mem[67],mem[66],mem[65],mem[64]} =32'b0000_0010_0100_00000_000_00010_0010011 ;
            {mem[71],mem[70],mem[69],mem[68]} =32'b0100001_00010_00000_010_00000_0100011 ;//sw

            {mem[75],mem[74],mem[73],mem[72]} =32'b0000_0100_0101_00000_000_00010_0010011 ;
            {mem[79],mem[78],mem[77],mem[76]} =32'b0100001_00010_00000_010_00100_0100011 ;//sw

            //////////////////////////////////////////////////////////////////////
            //x1 = max = 0
            {mem[83],mem[82],mem[81],mem[80]} =32'b0000_0000_0000_00000_000_00001_0010011 ; 
            // x2 = 10 (number of iterations)
            {mem[87],mem[86],mem[85],mem[84]} =32'b0000_0010_1000_00000_000_00010_0010011 ; 
            // x3 = i = 0
            {mem[91],mem[90],mem[89],mem[88]} =32'b0000_0000_0000_00000_000_00011_0010011 ; 
            // if i == 10, exit loop //beq x3, x2, end
            {mem[95],mem[94],mem[93],mem[92]} =32'b0000001_00011_00010_000_11110_1100011 ; 
            // x4 = array[i]
            {mem[99],mem[98],mem[97],mem[96]} =32'b0100000_00000_00011_010_00100_0000011 ;//lw
            //bge x4, x1, update_max // if array[i] >= max, update max
            {mem[103],mem[102],mem[101],mem[100]} =32'b0000000_00001_00100_101_01100_1100011 ; 
            // addi x3, x3, 4    // i++
            {mem[107],mem[106],mem[105],mem[104]} =32'b0000_0000_0100_00011_000_00011_0010011 ;
            //jal  loop
            {mem[111],mem[110],mem[109],mem[108]} =32'b1_1111111000_1_11111111_01111_1101111 ;


            //update_max:
            //addi x1, x4 , 0   // max = array[i]
            {mem[115],mem[114],mem[113],mem[112]} =32'b0000_0000_0000_00100_000_00001_0010011 ;
            // addi x3, x3, 4    // i++
            {mem[119],mem[118],mem[117],mem[116]} =32'b0000_0000_0100_00011_000_00011_0010011 ;
            //jal  loop
            {mem[123],mem[122],mem[121],mem[120]} =32'b1_1111110010_1_11111111_01111_1101111 ;
            // data_out <= {mem[3],mem[2],mem[1],mem[0]};
            

            //end LOOP
        end
    end
endmodule
